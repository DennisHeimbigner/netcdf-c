[0] /
[1] /.nczarr : (0) ||
