netcdf testmapnc4 {

group: _zarr {

  // group attributes:
  		:data = "" ;
  } // group _zarr
}
