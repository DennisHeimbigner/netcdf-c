[0] /testmapapi
[1] /testmapapi/.nczarr : (50) |7b0a22666f6f223a2034322c0a22626172223a20226170706c6573222c0a2262617a223a205b312c20322c20332c20345d7d|
[2] /testmapapi/data1 : (100) |000000000100000002000000030000000400000005000000060000000700000008000000090000000a0000000b0000000c0000000d0000000e0000000f000000100000001100000012000000130000001400000015000000160000001700000018000000|
[3] /testmapapi/meta1
[4] /testmapapi/meta1/.zarray : (34) |7b0a227368617065223a205b312c322c335d2c0a226474797065223a20223c31227d|
