./testmap.nzf
./testmap.nzf/.nczarr : ||
./testmap.nzf/meta1 : |{ "foo": 42, "bar": "apples", "baz": [1, 2, 3, 4]}|
