[1] /testmapapi/.nczarr : (0) ||
