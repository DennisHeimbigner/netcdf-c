./testmap.nzf
./testmap.nzf/meta2 : |{ "foo": 42, "bar": "apples", "baz": [1, 2, 3, 4], "extra": 137}|
./testmap.nzf/_nczarr : ||
./testmap.nzf/meta1 : |{ "foo": 42, "bar": "apples", "baz": [1, 2, 3, 4]}|
