netcdf ref_oldformat {
dimensions:
	lat = 8 ;
	_Anonymous_Dim_8 = 8 ;
	_Anonymous_Dim_10 = 10 ;
variables:
	int lat(_Anonymous_Dim_8) ;
		lat:_FillValue = -1 ;
		string lat:lat_attr = "latitude" ;
data:

 lat = 1, 2, 3, 4, 5, 6, 7, 8 ;

group: g1 {
  variables:
  	int pos(_Anonymous_Dim_8, _Anonymous_Dim_10) ;
  		pos:_FillValue = -1 ;
  		string pos:pos_attr = "latXlon" ;

  // group attributes:
  		:g1_attr = 17 ;
  data:

   pos =
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _,
  _, _, _, _, _, _, _, _, _, _ ;
  } // group g1
}
