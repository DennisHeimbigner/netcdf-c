./testmap.nzf
./testmap.nzf/_nczarr : ||
