netcdf testnc4 {
}
