netcdf testnc4 {
dimensions:
	meta1 = UNLIMITED ; // (50 currently)
	meta2 = UNLIMITED ; // (64 currently)
variables:
	ubyte meta1(meta1) ;
		meta1:_FillValue = 0UB ;
		meta1:text = "{\n\"foo\": 42,\n\"bar\": \"apples\",\n\"baz\": [1, 2, 3, 4]}" ;
	ubyte meta2(meta2) ;
		meta2:_FillValue = 0UB ;
		meta2:text = "{\n\"foo\": 42,\n\"bar\": \"apples\",\n\"baz\": [1, 2, 3, 4],\n\"extra\": 137}" ;
data:

 meta1 = 123, 10, 34, 102, 111, 111, 34, 58, 32, 52, 50, 44, 10, 34, 98, 97, 
    114, 34, 58, 32, 34, 97, 112, 112, 108, 101, 115, 34, 44, 10, 34, 98, 97, 
    122, 34, 58, 32, 91, 49, 44, 32, 50, 44, 32, 51, 44, 32, 52, 93, 125 ;

 meta2 = 123, 10, 34, 102, 111, 111, 34, 58, 32, 52, 50, 44, 10, 34, 98, 97, 
    114, 34, 58, 32, 34, 97, 112, 112, 108, 101, 115, 34, 44, 10, 34, 98, 97, 
    122, 34, 58, 32, 91, 49, 44, 32, 50, 44, 32, 51, 44, 32, 52, 93, 44, 10, 
    34, 101, 120, 116, 114, 97, 34, 58, 32, 49, 51, 55, 125 ;
}
