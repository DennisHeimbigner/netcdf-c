[0] /testmapapi
[1] /testmapapi/.nczarr : (50) |7b0a22666f6f223a2034322c0a22626172223a20226170706c6573222c0a2262617a223a205b312c20322c20332c20345d7d|
[2] /testmapapi/meta1
[3] /testmapapi/meta1/.zarray : (34) |7b0a227368617065223a205b312c322c335d2c0a226474797065223a20223c31227d|
