netcdf testmap {

group: _nczarr {
  } // group _nczarr

group: meta1 {

  group: _zarray {

    // group attributes:
    		:data = "{\n\"foo\": 42,\n\"bar\": \"apples\",\n\"baz\": [1, 2, 3, 4]}" ;
    } // group _zarray
  } // group meta1

group: meta2 {

  group: _nczvar {

    // group attributes:
    		:data = "{\n\"foo\": 42,\n\"bar\": \"apples\",\n\"baz\": [1, 2, 3, 4],\n\"extra\": 137}" ;
    } // group _nczvar
  } // group meta2
}
