netcdf testmapnc4 {

group: _nczarr {

  // group attributes:
  		:data = "" ;
  } // group _nczarr
}
