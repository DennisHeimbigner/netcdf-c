[0] /testmapapi
[1] /testmapapi/.nczarr : (0) ||
