[1] / : (0) ||
[0] /.nczarr : (0) ||
