[1] /testmapapi/.nczarr : (50) |{
"foo": 42,
"bar": "apples",
"baz": [1, 2, 3, 4]}|
[2] /testmapapi/data1 : (100) |000000000100000002000000030000000400000005000000060000000700000008000000090000000a0000000b0000000c0000000d0000000e0000000f000000100000001100000012000000130000001400000015000000160000001700000018000000|
[4] /testmapapi/meta1/.zarray : (34) |{
"shape": [1,2,3],
"dtype": "<1"}|
